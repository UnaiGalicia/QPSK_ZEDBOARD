--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   07:23:48 01/07/2014
-- Design Name:   
-- Module Name:   C:/Users/hamster/Projects/FPGA/egokitu_test/egokitu_tb.vhd
-- Project Name:  egokitu_test
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: egokitu_test
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types- always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY egokitu_tb IS
END egokitu_tb;
 
ARCHITECTURE behavior OF egokitu_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
	COMPONENT qpsk_egokitu
	PORT(
		   audio_serie : in STD_LOGIC_VECTOR (31 downto 0);
           audio_L : out STD_LOGIC_VECTOR (23 downto 0);
           audio_R : out STD_LOGIC_VECTOR (23 downto 0);
           nsample: in STD_LOGIC;
           axi_tvalid: in STD_LOGIC;
           axi_tready: out STD_LOGIC;
           clk : in STD_LOGIC
           
		);
	END COMPONENT;    

   --Inputs
   signal clk : std_logic := '0';
   signal audio_serie : std_logic_vector (31 downto 0);
   signal nsample : std_logic;
   signal axi_tvalid : std_logic;
   --signal AC_GPIO1 : std_logic := '0';

	--BiDirs
   --signal AC_SDA : std_logic;

 	--Outputs
   signal	audio_L	:	std_logic_vector(23 downto 0);
   signal	audio_R	:	std_logic_vector(23 downto 0);
   signal	axi_tready	:	std_logic;
   
 

   --signal lr_stim  : std_logic_vector(63 downto 0) := x"FFFFFFFF00000000";
   --signal d_stim   : std_logic_vector(63 downto 0) := x"4000000040000000";
   -- Clock period definitions
   --constant clk_period : time := 10 ns;
   constant	clk48_period : time := 20 ns;
BEGIN
   --AC_SDA <= 'H';
   
	-- Instantiate the Unit Under Test (UUT)
   uut: qpsk_egokitu PORT MAP (
		  audio_serie => audio_serie,
          audio_L => audio_L,
          audio_R => audio_R,
          nsample => nsample,
          axi_tvalid => axi_tvalid,
          axi_tready => axi_tready,
          clk => clk
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk48_period/2;
		clk <= '1';
		wait for clk48_period/2;
   end process;
 
   --AC_GPIO3 <= lr_stim(lr_stim'high);
   --AC_GPIO1 <= d_stim(d_stim'high);


-- simulate the clocks generated by the codec chip.   
 simulazioa : process
   begin
   
	nsample <= '0';
	axi_tvalid <='0';
	audio_serie <= "00000000000000010000000000000011";
	wait for 60 ns;
	
	nsample <= '1';
	axi_tvalid <='0';
	audio_serie <= "00000000000000010000000000000011";
	wait for 60 ns;
	
    nsample <= '0';
	axi_tvalid <='0';
	audio_serie <= "00000000000000010000000000000011";
	wait for 60 ns;
	
	nsample <= '0';
	axi_tvalid <='1';
	audio_serie <= "00000000000001110000000011000011";
	wait for 60 ns;
	
	nsample <= '0';
	axi_tvalid <='0';
	audio_serie <= "00000000000000010000000000000011";
	wait for 60 ns;
	
	nsample <= '1';
	axi_tvalid <='0';
	audio_serie <= "00000000101111110110000011000011";
	wait for 60 ns;
	
	nsample <= '0';
	axi_tvalid <='1';
	audio_serie <= "00000000101111110110000011000011";
	wait for 60 ns;
	
	nsample <= '0';
	axi_tvalid <='0';
	audio_serie <= "00000000101111110110000011000011";
	wait for 60 ns;
	
   end process;
   -- Stimulus process
   stim_proc: process
   begin		
      wait;
   end process;

END;
